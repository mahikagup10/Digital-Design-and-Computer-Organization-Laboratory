module testbench;

reg clk, reset;

endmodule